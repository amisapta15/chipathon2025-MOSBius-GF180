** sch_path: /foss/designs/Chipathon2025_gf180/gf180_examples/RO/xschem/3_stage_RO_tb_tran.sch
**.subckt 3_stage_RO_tb_tran
x1 VDD VSS n1 3_stage_RO
V1 VSS GND 0
V2 VDD VSS 3.3
* noconn n1
**** begin user architecture code

.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/smbb000149.ngspice typical



.tran 1n 10u
.save all
.ic V(n1)=0


**** end user architecture code
**.ends

* expanding   symbol:  3_stage_RO.sym # of pins=3
** sym_path: /foss/designs/Chipathon2025_gf180/gf180_examples/RO/xschem/3_stage_RO.sym
** sch_path: /foss/designs/Chipathon2025_gf180/gf180_examples/RO/xschem/3_stage_RO.sch
.subckt 3_stage_RO VDD VSS n1
*.iopin VDD
*.iopin VSS
*.iopin n1
x1 n1 VDD VSS n2 inverter
x2 n2 VDD VSS n3 inverter
x3 n3 VDD VSS n1 inverter
.ends


* expanding   symbol:  /foss/designs/Chipathon2025_gf180/gf180_examples/inverter/xschem/inverter.sym # of pins=4
** sym_path: /foss/designs/Chipathon2025_gf180/gf180_examples/inverter/xschem/inverter.sym
** sch_path: /foss/designs/Chipathon2025_gf180/gf180_examples/inverter/xschem/inverter.sch
.subckt inverter Vin VDD VSS Vout
*.ipin Vin
*.iopin VDD
*.iopin VSS
*.iopin Vout
XM1 Vout Vin VSS VSS nfet_03v3 L=1u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 Vout Vin VDD VDD pfet_03v3 L=1u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
