* Extracted by KLayout with GF180MCU LVS runset on : 04/09/2025 22:03

.SUBCKT 3_stage_RO VSS n1 VDD
M$1 \$2 n1 VDD VDD pfet_03v3 L=1U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$2 \$3 \$2 VDD VDD pfet_03v3 L=1U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$3 n1 \$3 VDD VDD pfet_03v3 L=1U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$4 \$2 n1 VSS VSS nfet_03v3 L=1U W=3U AS=1.83P AD=1.83P PS=7.22U PD=7.22U
M$5 \$3 \$2 VSS VSS nfet_03v3 L=1U W=3U AS=1.83P AD=1.83P PS=7.22U PD=7.22U
M$6 n1 \$3 VSS VSS nfet_03v3 L=1U W=3U AS=1.83P AD=1.83P PS=7.22U PD=7.22U
.ENDS 3_stage_RO
